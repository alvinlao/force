library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity sad is
	generic(
		pixel_buffer_base : std_logic_vector := x"00000000";
		win_size_x: integer := 20;
		win_size_y: integer := 20;
		block_size_x: integer := 7;
		block_size_y: integer := 7;
		step_x: integer := 1;
		step_y: integer := 1		
	);	
	port (
		clk		: in std_logic;
		reset_n	: in std_logic;
		
		start 	: in std_logic;
		ready 	: out std_logic;
		
		posX 	: out std_logic_vector(8 downto 0);
		posY 	: out std_logic_vector(7 downto 0);
		acc		: out std_logic_vector(15 downto 0);
				
		master_addr : out std_logic_vector(31 downto 0);
		master_rd_en : out std_logic;
		master_wr_en : out std_logic;
		master_be : out std_logic_vector(1 downto 0);
		master_readdata : in std_logic_vector(15 downto 0);
		master_writedata: out  std_logic_vector(15 downto 0);
		master_waitrequest : in std_logic
	);
end sad;

architecture bhv of sad is
	constant SCREEN_WIDTH 	: integer := 320;
	constant SCREEN_HEIGHT 	: integer := 240;
	constant SAD_SIZE 		: integer := 65536;
	
	type StatesType				is (Standby,Loading,CalculatingSAD, AddingSAD,Picking);
	type WindowType 			is array (0 to win_size_x, 0 to win_size_y) of std_logic_vector(15 downto 0);
	type BlockType 				is array (0 to block_size_x, 0 to block_size_y) of std_logic_vector(15 downto 0);
	type SadBlockType 			is array (0 to block_size_x-1, 0 to block_size_y-1) of integer range 0 to SAD_SIZE;
	type SadWindowType 			is array (0 to ((win_size_x - block_size_x)/step_x), 0 to (win_size_y - block_size_y)/step_y) of SadBlockType;
	type SADForEachBlocksType	is array (0 to ((win_size_x - block_size_x)/step_x), 0 to (win_size_y - block_size_y)/step_y) of integer range 0 to SAD_SIZE;
	
    signal current_state 	: StatesType := Standby;
	signal next_state 		: StatesType := Standby;
	
	signal Window 			: WindowType;
	
	signal windowStartX 	: integer range 0 to (SCREEN_WIDTH - win_size_x);
	signal windowStartY 	: integer range 0 to (SCREEN_HEIGHT - win_size_y);
	
	signal ReferenceBlock 	: BlockType;
	signal SADForEachBlock 	: SADForEachBlocksType;	
	signal SADCollection 	: SadWindowType;
	
	begin
	  
	process (clk, reset_n)

	variable nextX : integer range 0 to SCREEN_WIDTH;
		variable nextY : integer range 0 to SCREEN_HEIGHT;
		variable candidateRow : integer range 0 to ((win_size_x - block_size_x)/step_x);
		variable candidateCol : integer range 0 to ((win_size_y - block_size_y)/step_y);
		variable candidateSAD : integer range 0 to SAD_SIZE := SAD_SIZE;
		variable load_waiting : std_logic;

	begin
		if (reset_n = '0') then
			current_state <= Standby;
			next_state <= Standby;
			ready <= '0';
		elsif rising_edge(clk) then
			next_state <= current_state;
			master_wr_en <= '0';
			master_rd_en <= '0';
						
			case (current_state) is
				when Standby => 
						if (start = '1') then
							next_state <= Loading;
							nextX := 0;
							nextY := 0;
							load_waiting := '0';
							ready <= '0';
						end if;

				when Loading =>
					ready <= '0';
					if (load_waiting = '1') then
						if (master_waitrequest = '0') then
							load_waiting := '0';
							master_wr_en <= '0';
							master_rd_en <= '0';

							Window(nextX,nextY) <= master_readdata;
							
							nextX := nextX+1;
							if(nextX = block_size_x) then
								nextX := 0;
								nextY := nextY +1;
								
								if (nextY = block_size_y) then
									next_state <= CalculatingSAD;
									load_waiting := '1';
								end if;
							end if;
						else
							master_addr <= std_logic_vector(unsigned(pixel_buffer_base) + unsigned(to_unsigned(windowStartX + nextX, 9)) & unsigned(to_unsigned(windowStartY + nextY, 8)) & '0');	
							master_be <= "11";  -- byte enable
							master_wr_en <= '0';
							master_rd_en <= '1';
						end if;
					else
						master_addr <= std_logic_vector(unsigned(pixel_buffer_base) + unsigned(to_unsigned(windowStartX + nextX, 9)) & unsigned(to_unsigned(windowStartY + nextY, 8)) & '0');	
						master_be <= "11";  -- byte enable
						master_wr_en <= '0';
						master_rd_en <= '1';
						
						load_waiting := '1';
					end if;
		
				when CalculatingSAD =>
					ready <= '0';
					
					for WIN_ROW in 0 to ((win_size_x - block_size_x)/step_x) loop
						for WIN_COL in 0 to ((win_size_y - block_size_y)/step_y) loop
							for BLK_ROW in 0 to (block_size_x-1) loop
								for BLK_COL in 0 to (block_size_y-1) loop
									SADCollection(WIN_ROW,WIN_COL)(BLK_ROW,BLK_COL) <= to_integer(
										(unsigned((signed('0'&Window((WIN_ROW*step_x)+BLK_ROW,(WIN_COL*step_y)+BLK_COL)(15 downto 11)) - signed('0'&ReferenceBlock(WIN_ROW+BLK_ROW,WIN_COL+BLK_COL)(15 downto 11)))) and B"01_1111") + 
										(unsigned((signed('0'&Window((WIN_ROW*step_x)+BLK_ROW,(WIN_COL*step_y)+BLK_COL)(10 downto 5)) - signed('0'&ReferenceBlock(WIN_ROW+BLK_ROW,WIN_COL+BLK_COL)(10 downto 5)))) and B"011_1111" ) + 
										(unsigned((signed('0'&Window((WIN_ROW*step_x)+BLK_ROW,(WIN_COL*step_y)+BLK_COL)(4 downto 0)) - signed('0'&ReferenceBlock(WIN_ROW+BLK_ROW,WIN_COL+BLK_COL)(4 downto 0)))) and B"01_1111")
										);
								end loop;																
							end loop;													
						end loop;						
					end loop;
					
					nextX := 0;
					nextY := 0;
					next_state <= AddingSAD;
					
				when AddingSAD =>
					ready <= '0';
				
					for WIN_ROW in 0 to ((win_size_x - block_size_x)/step_x) loop
						for WIN_COL in 0 to ((win_size_y - block_size_y)/step_y) loop
						
							SADForEachBlock(WIN_ROW,WIN_COL) <= SADForEachBlock(WIN_ROW,WIN_COL) + SADCollection(WIN_ROW,WIN_COL)(nextX,nextY);
							
						end loop;						
					end loop;
					
					nextX := nextX+1;
					if(nextX = block_size_x) then
						nextX := 0;
						nextY := nextY +1;
						
						if (nextY = block_size_y) then
							candidateSAD := SAD_SIZE;
							next_state <= Picking;
						end if;
					end if;
					
				when Picking =>
					
					for WIN_ROW in 0 to ((win_size_x - block_size_x)/step_x) loop
						for WIN_COL in 0 to ((win_size_y - block_size_y)/step_y) loop
						
							if (SADForEachBlock(WIN_ROW,WIN_COL) < candidateSAD) then
								candidateSAD := SADForEachBlock(WIN_ROW,WIN_COL);
								candidateRow := WIN_ROW;
								candidateCol := WIN_COL;
							end if;
							
						end loop;						
					end loop;

					posX <= std_logic_vector(to_unsigned((candidateRow*step_x)+(block_size_x/2),9));
					posY <= std_logic_vector(to_unsigned((candidateCol*step_y)+(block_size_y/2),8));
					acc <= std_logic_vector(to_unsigned(candidateSAD,16));
					ready <= '1';
					next_state <= Standby;
					
				when others=>
					-- why are we here?
					next_state <= Standby;
			end case;
		end if;	
	end process;	
				
end bhv;
